/* 19_vector5.v
 * aaaaa_bbbbb_ccccc_ddddd_eeeee
 * abcde_abcde_abcde_abcde_abcde
 * bit24 --> bit0
 */

module top_module (
    input a, b, c, d, e,
    output [24:0] out );//

    // The output is XNOR of two vectors created by 
    // concatenating and replicating the five inputs.
    // assign out = ~{ ... } ^ { ... };
    assign out = ~{ {5{a}},{5{b}},{5{c}},{5{d}},{5{e}} } ^ { 5{a,b,c,d,e} };

	// wire [24:0] top, bottom;
	// assign top    = { {5{a}}, {5{b}}, {5{c}}, {5{d}}, {5{e}} };
	// assign bottom = {5{a,b,c,d,e}};
	// assign out = ~top ^ bottom;	// Bitwise XNOR

endmodule
